LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;	
ENTITY Finaladder IS
  PORT (
  		clk			: IN 		STD_LOGIC;
		adder			: IN		STD_LOGIC_VECTOR(31 DOWNTO 0);
		multiply		: IN		STD_LOGIC_VECTOR(31 DOWNTO 0)

);		
END ENTITY Finaladder;


ARCHITECTURE structure OF Finaladder IS

BEGIN

END;