
module uart (
	reset_reset_n);	

	input		reset_reset_n;
endmodule
